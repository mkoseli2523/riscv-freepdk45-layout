/home/mkoseli2/Desktop/ece425.work/release/mp_pnr/provided/stdcells.lef